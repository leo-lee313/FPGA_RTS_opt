// megafunction wizard: %LPM_MUX%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_MUX 

// ============================================================
// File Name: muxer7.v
// Megafunction Name(s):
// 			LPM_MUX
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.0.1 Build 232 06/12/2013 SP 1 SJ Full Version
// ************************************************************

//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module muxer7 (
	clock,
	data0x,
	data1x,
	data2x,
	data3x,
	data4x,
	data5x,
	data6x,
	data7x,
	sel,
	result);

	input	  clock;
	input	[63:0]  data0x;
	input	[63:0]  data1x;
	input	[63:0]  data2x;
	input	[63:0]  data3x;
	input	[63:0]  data4x;
	input	[63:0]  data5x;
	input	[63:0]  data6x;
	input	[63:0]  data7x;
	input	[2:0]  sel;
	output	[63:0]  result;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix V"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "1"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "1"
// Retrieval info: CONSTANT: LPM_SIZE NUMERIC "8"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "64"
// Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "3"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: data0x 0 0 64 0 INPUT NODEFVAL "data0x[63..0]"
// Retrieval info: USED_PORT: data1x 0 0 64 0 INPUT NODEFVAL "data1x[63..0]"
// Retrieval info: USED_PORT: data2x 0 0 64 0 INPUT NODEFVAL "data2x[63..0]"
// Retrieval info: USED_PORT: data3x 0 0 64 0 INPUT NODEFVAL "data3x[63..0]"
// Retrieval info: USED_PORT: data4x 0 0 64 0 INPUT NODEFVAL "data4x[63..0]"
// Retrieval info: USED_PORT: data5x 0 0 64 0 INPUT NODEFVAL "data5x[63..0]"
// Retrieval info: USED_PORT: data6x 0 0 64 0 INPUT NODEFVAL "data6x[63..0]"
// Retrieval info: USED_PORT: data7x 0 0 64 0 INPUT NODEFVAL "data7x[63..0]"
// Retrieval info: USED_PORT: result 0 0 64 0 OUTPUT NODEFVAL "result[63..0]"
// Retrieval info: USED_PORT: sel 0 0 3 0 INPUT NODEFVAL "sel[2..0]"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 64 0 data0x 0 0 64 0
// Retrieval info: CONNECT: @data 0 0 64 64 data1x 0 0 64 0
// Retrieval info: CONNECT: @data 0 0 64 128 data2x 0 0 64 0
// Retrieval info: CONNECT: @data 0 0 64 192 data3x 0 0 64 0
// Retrieval info: CONNECT: @data 0 0 64 256 data4x 0 0 64 0
// Retrieval info: CONNECT: @data 0 0 64 320 data5x 0 0 64 0
// Retrieval info: CONNECT: @data 0 0 64 384 data6x 0 0 64 0
// Retrieval info: CONNECT: @data 0 0 64 448 data7x 0 0 64 0
// Retrieval info: CONNECT: @sel 0 0 3 0 sel 0 0 3 0
// Retrieval info: CONNECT: result 0 0 64 0 @result 0 0 64 0
// Retrieval info: GEN_FILE: TYPE_NORMAL muxer7.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL muxer7.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL muxer7.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL muxer7.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL muxer7_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL muxer7_bb.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL muxer7_syn.v TRUE
// Retrieval info: LIB_FILE: lpm
